//NOTE: This is based on this:
// https://github.com/algofoogle/raybox/blob/main/src/rtl/lzc_b.v
//...in this case, hard-coded for 24-bit inputs, i.e. Q12.12.

`default_nettype none
`timescale 1ns / 1ps


module lzc(
  input [23:0] i_data,
  output [4:0] o_lzc      // 0..24 is normal.
);

  function [4:0] f_lzc(input [23:0] data);
    casez (i_data)
      24'b1???????????????????????:  f_lzc =  0;
      24'b01??????????????????????:  f_lzc =  1;
      24'b001?????????????????????:  f_lzc =  2;
      24'b0001????????????????????:  f_lzc =  3;
      24'b00001???????????????????:  f_lzc =  4;
      24'b000001??????????????????:  f_lzc =  5;
      24'b0000001?????????????????:  f_lzc =  6;
      24'b00000001????????????????:  f_lzc =  7;
      24'b000000001???????????????:  f_lzc =  8;
      24'b0000000001??????????????:  f_lzc =  9;
      24'b00000000001?????????????:  f_lzc = 10;
      24'b000000000001????????????:  f_lzc = 11;
      24'b0000000000001???????????:  f_lzc = 12;
      24'b00000000000001??????????:  f_lzc = 13;
      24'b000000000000001?????????:  f_lzc = 14;
      24'b0000000000000001????????:  f_lzc = 15;
      24'b00000000000000001???????:  f_lzc = 16;
      24'b000000000000000001??????:  f_lzc = 17;
      24'b0000000000000000001?????:  f_lzc = 18;
      24'b00000000000000000001????:  f_lzc = 19;
      24'b000000000000000000001???:  f_lzc = 20;
      24'b0000000000000000000001??:  f_lzc = 21;
      24'b00000000000000000000001?:  f_lzc = 22;
      24'b000000000000000000000001:  f_lzc = 23;
      24'b000000000000000000000000:  f_lzc = 24;
    endcase

  endfunction

  assign o_lzc = f_lzc(i_data);

endmodule
