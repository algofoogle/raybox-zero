//NOTE: This is based on this:
// https://github.com/algofoogle/raybox/blob/main/src/rtl/lzc_b.v
//...in this case, hard-coded for 20-bit inputs, i.e. Q10.10.

`default_nettype none
`timescale 1ns / 1ps

`include "fixed_point_params.v"

`define INRANGE [`Qm-1:-`Qn]

module lzc(
  input `INRANGE i_data,
  output [4:0] o_lzc      // 0..20 is normal.
);

  function [4:0] f_lzc(input `INRANGE data);
    casez (i_data)
      //SMELL: This is probably a sloppy way to do this, and it is currently hard-coded for 20-bit inputs only:
      20'b1???????????????????:  f_lzc =  0;
      20'b01??????????????????:  f_lzc =  1;
      20'b001?????????????????:  f_lzc =  2;
      20'b0001????????????????:  f_lzc =  3;
      20'b00001???????????????:  f_lzc =  4;
      20'b000001??????????????:  f_lzc =  5;
      20'b0000001?????????????:  f_lzc =  6;
      20'b00000001????????????:  f_lzc =  7;
      20'b000000001???????????:  f_lzc =  8;
      20'b0000000001??????????:  f_lzc =  9;
      20'b00000000001?????????:  f_lzc = 10;
      20'b000000000001????????:  f_lzc = 11;
      20'b0000000000001???????:  f_lzc = 12;
      20'b00000000000001??????:  f_lzc = 13;
      20'b000000000000001?????:  f_lzc = 14;
      20'b0000000000000001????:  f_lzc = 15;
      20'b00000000000000001???:  f_lzc = 16;
      20'b000000000000000001??:  f_lzc = 17;
      20'b0000000000000000001?:  f_lzc = 18;
      20'b00000000000000000001:  f_lzc = 19;
      20'b00000000000000000000:  f_lzc = 20;
    endcase

  endfunction

  assign o_lzc = f_lzc(i_data);

endmodule
